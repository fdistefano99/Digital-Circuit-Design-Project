
    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end projecttb;